// DE10_Standard_VIP_Qsys.v

// Generated using ACDS version 16.1 200

`timescale 1 ps / 1 ps
module DE10_Standard_VIP_Qsys (
		input  wire        alt_vip_cl_cvi_0_clocked_video_vid_clk,            // alt_vip_cl_cvi_0_clocked_video.vid_clk
		input  wire [7:0]  alt_vip_cl_cvi_0_clocked_video_vid_data,           //                               .vid_data
		input  wire        alt_vip_cl_cvi_0_clocked_video_vid_de,             //                               .vid_de
		input  wire        alt_vip_cl_cvi_0_clocked_video_vid_datavalid,      //                               .vid_datavalid
		input  wire        alt_vip_cl_cvi_0_clocked_video_vid_locked,         //                               .vid_locked
		input  wire        alt_vip_cl_cvi_0_clocked_video_vid_f,              //                               .vid_f
		input  wire        alt_vip_cl_cvi_0_clocked_video_vid_v_sync,         //                               .vid_v_sync
		input  wire        alt_vip_cl_cvi_0_clocked_video_vid_h_sync,         //                               .vid_h_sync
		input  wire [7:0]  alt_vip_cl_cvi_0_clocked_video_vid_color_encoding, //                               .vid_color_encoding
		input  wire [7:0]  alt_vip_cl_cvi_0_clocked_video_vid_bit_width,      //                               .vid_bit_width
		output wire        alt_vip_cl_cvi_0_clocked_video_sof,                //                               .sof
		output wire        alt_vip_cl_cvi_0_clocked_video_sof_locked,         //                               .sof_locked
		output wire        alt_vip_cl_cvi_0_clocked_video_refclk_div,         //                               .refclk_div
		output wire        alt_vip_cl_cvi_0_clocked_video_clipping,           //                               .clipping
		output wire        alt_vip_cl_cvi_0_clocked_video_padding,            //                               .padding
		output wire        alt_vip_cl_cvi_0_clocked_video_overflow,           //                               .overflow
		input  wire        alt_vip_itc_0_clocked_video_vid_clk,               //    alt_vip_itc_0_clocked_video.vid_clk
		output wire [23:0] alt_vip_itc_0_clocked_video_vid_data,              //                               .vid_data
		output wire        alt_vip_itc_0_clocked_video_underflow,             //                               .underflow
		output wire        alt_vip_itc_0_clocked_video_vid_datavalid,         //                               .vid_datavalid
		output wire        alt_vip_itc_0_clocked_video_vid_v_sync,            //                               .vid_v_sync
		output wire        alt_vip_itc_0_clocked_video_vid_h_sync,            //                               .vid_h_sync
		output wire        alt_vip_itc_0_clocked_video_vid_f,                 //                               .vid_f
		output wire        alt_vip_itc_0_clocked_video_vid_h,                 //                               .vid_h
		output wire        alt_vip_itc_0_clocked_video_vid_v,                 //                               .vid_v
		input  wire        clk_clk,                                           //                            clk.clk
		output wire        clk_aud_clk,                                       //                        clk_aud.clk
		output wire        clk_sdram_clk,                                     //                      clk_sdram.clk
		output wire        clk_vga_clk,                                       //                        clk_vga.clk
		input  wire        reset_reset_n,                                     //                          reset.reset_n
		output wire [12:0] sdram_wire_addr,                                   //                     sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                                     //                               .ba
		output wire        sdram_wire_cas_n,                                  //                               .cas_n
		output wire        sdram_wire_cke,                                    //                               .cke
		output wire        sdram_wire_cs_n,                                   //                               .cs_n
		inout  wire [15:0] sdram_wire_dq,                                     //                               .dq
		output wire [1:0]  sdram_wire_dqm,                                    //                               .dqm
		output wire        sdram_wire_ras_n,                                  //                               .ras_n
		output wire        sdram_wire_we_n                                    //                               .we_n
	);

	wire         alt_vip_cl_vfb_0_dout_valid;                  // alt_vip_cl_vfb_0:dout_valid -> alt_vip_cl_crs_0:din_valid
	wire  [15:0] alt_vip_cl_vfb_0_dout_data;                   // alt_vip_cl_vfb_0:dout_data -> alt_vip_cl_crs_0:din_data
	wire         alt_vip_cl_vfb_0_dout_ready;                  // alt_vip_cl_crs_0:din_ready -> alt_vip_cl_vfb_0:dout_ready
	wire         alt_vip_cl_vfb_0_dout_startofpacket;          // alt_vip_cl_vfb_0:dout_startofpacket -> alt_vip_cl_crs_0:din_startofpacket
	wire         alt_vip_cl_vfb_0_dout_endofpacket;            // alt_vip_cl_vfb_0:dout_endofpacket -> alt_vip_cl_crs_0:din_endofpacket
	wire         alt_vip_cl_crs_0_dout_valid;                  // alt_vip_cl_crs_0:dout_valid -> alt_vip_cl_csc_0:din_valid
	wire  [23:0] alt_vip_cl_crs_0_dout_data;                   // alt_vip_cl_crs_0:dout_data -> alt_vip_cl_csc_0:din_data
	wire         alt_vip_cl_crs_0_dout_ready;                  // alt_vip_cl_csc_0:din_ready -> alt_vip_cl_crs_0:dout_ready
	wire         alt_vip_cl_crs_0_dout_startofpacket;          // alt_vip_cl_crs_0:dout_startofpacket -> alt_vip_cl_csc_0:din_startofpacket
	wire         alt_vip_cl_crs_0_dout_endofpacket;            // alt_vip_cl_crs_0:dout_endofpacket -> alt_vip_cl_csc_0:din_endofpacket
	wire         alt_vip_clip_1_dout_valid;                    // alt_vip_clip_1:dout_valid -> alt_vip_cl_vfb_0:din_valid
	wire  [15:0] alt_vip_clip_1_dout_data;                     // alt_vip_clip_1:dout_data -> alt_vip_cl_vfb_0:din_data
	wire         alt_vip_clip_1_dout_ready;                    // alt_vip_cl_vfb_0:din_ready -> alt_vip_clip_1:dout_ready
	wire         alt_vip_clip_1_dout_startofpacket;            // alt_vip_clip_1:dout_startofpacket -> alt_vip_cl_vfb_0:din_startofpacket
	wire         alt_vip_clip_1_dout_endofpacket;              // alt_vip_clip_1:dout_endofpacket -> alt_vip_cl_vfb_0:din_endofpacket
	wire         alt_vip_cl_dil_0_dout_valid;                  // alt_vip_cl_dil_0:dout_valid -> alt_vip_clip_1:din_valid
	wire  [15:0] alt_vip_cl_dil_0_dout_data;                   // alt_vip_cl_dil_0:dout_data -> alt_vip_clip_1:din_data
	wire         alt_vip_cl_dil_0_dout_ready;                  // alt_vip_clip_1:din_ready -> alt_vip_cl_dil_0:dout_ready
	wire         alt_vip_cl_dil_0_dout_startofpacket;          // alt_vip_cl_dil_0:dout_startofpacket -> alt_vip_clip_1:din_startofpacket
	wire         alt_vip_cl_dil_0_dout_endofpacket;            // alt_vip_cl_dil_0:dout_endofpacket -> alt_vip_clip_1:din_endofpacket
	wire         alt_vip_cl_csc_0_dout_valid;                  // alt_vip_cl_csc_0:dout_valid -> alt_vip_scl_0:din_valid
	wire  [23:0] alt_vip_cl_csc_0_dout_data;                   // alt_vip_cl_csc_0:dout_data -> alt_vip_scl_0:din_data
	wire         alt_vip_cl_csc_0_dout_ready;                  // alt_vip_scl_0:din_ready -> alt_vip_cl_csc_0:dout_ready
	wire         alt_vip_cl_csc_0_dout_startofpacket;          // alt_vip_cl_csc_0:dout_startofpacket -> alt_vip_scl_0:din_startofpacket
	wire         alt_vip_cl_csc_0_dout_endofpacket;            // alt_vip_cl_csc_0:dout_endofpacket -> alt_vip_scl_0:din_endofpacket
	wire         alt_vip_scl_0_dout_valid;                     // alt_vip_scl_0:dout_valid -> alt_vip_itc_0:is_valid
	wire  [23:0] alt_vip_scl_0_dout_data;                      // alt_vip_scl_0:dout_data -> alt_vip_itc_0:is_data
	wire         alt_vip_scl_0_dout_ready;                     // alt_vip_itc_0:is_ready -> alt_vip_scl_0:dout_ready
	wire         alt_vip_scl_0_dout_startofpacket;             // alt_vip_scl_0:dout_startofpacket -> alt_vip_itc_0:is_sop
	wire         alt_vip_scl_0_dout_endofpacket;               // alt_vip_scl_0:dout_endofpacket -> alt_vip_itc_0:is_eop
	wire         alt_vip_cl_cps_0_dout_0_valid;                // alt_vip_cl_cps_0:dout_0_valid -> alt_vip_cl_dil_0:din_valid
	wire  [15:0] alt_vip_cl_cps_0_dout_0_data;                 // alt_vip_cl_cps_0:dout_0_data -> alt_vip_cl_dil_0:din_data
	wire         alt_vip_cl_cps_0_dout_0_ready;                // alt_vip_cl_dil_0:din_ready -> alt_vip_cl_cps_0:dout_0_ready
	wire         alt_vip_cl_cps_0_dout_0_startofpacket;        // alt_vip_cl_cps_0:dout_0_startofpacket -> alt_vip_cl_dil_0:din_startofpacket
	wire         alt_vip_cl_cps_0_dout_0_endofpacket;          // alt_vip_cl_cps_0:dout_0_endofpacket -> alt_vip_cl_dil_0:din_endofpacket
	wire         alt_vip_cl_cvi_0_dout_0_valid;                // alt_vip_cl_cvi_0:dout_0_valid -> alt_vip_cl_cps_0:din_0_valid
	wire   [7:0] alt_vip_cl_cvi_0_dout_0_data;                 // alt_vip_cl_cvi_0:dout_0_data -> alt_vip_cl_cps_0:din_0_data
	wire         alt_vip_cl_cvi_0_dout_0_ready;                // alt_vip_cl_cps_0:din_0_ready -> alt_vip_cl_cvi_0:dout_0_ready
	wire         alt_vip_cl_cvi_0_dout_0_startofpacket;        // alt_vip_cl_cvi_0:dout_0_startofpacket -> alt_vip_cl_cps_0:din_0_startofpacket
	wire         alt_vip_cl_cvi_0_dout_0_endofpacket;          // alt_vip_cl_cvi_0:dout_0_endofpacket -> alt_vip_cl_cps_0:din_0_endofpacket
	wire         pll_0_outclk1_clk;                            // pll_0:outclk_1 -> [alt_vip_cl_cps_0:main_clock, alt_vip_cl_crs_0:main_clock, alt_vip_cl_csc_0:main_clock, alt_vip_cl_cvi_0:main_clock_clk, alt_vip_cl_dil_0:av_st_clock, alt_vip_cl_vfb_0:main_clock, alt_vip_cl_vfb_0:mem_clock, alt_vip_clip_1:main_clock, alt_vip_itc_0:is_clk, alt_vip_scl_0:main_clock, mm_interconnect_0:pll_0_outclk1_clk, rst_controller:clk, sdram:clk]
	wire         alt_vip_cl_vfb_0_mem_master_rd_waitrequest;   // mm_interconnect_0:alt_vip_cl_vfb_0_mem_master_rd_waitrequest -> alt_vip_cl_vfb_0:mem_master_rd_waitrequest
	wire  [31:0] alt_vip_cl_vfb_0_mem_master_rd_readdata;      // mm_interconnect_0:alt_vip_cl_vfb_0_mem_master_rd_readdata -> alt_vip_cl_vfb_0:mem_master_rd_readdata
	wire  [31:0] alt_vip_cl_vfb_0_mem_master_rd_address;       // alt_vip_cl_vfb_0:mem_master_rd_address -> mm_interconnect_0:alt_vip_cl_vfb_0_mem_master_rd_address
	wire         alt_vip_cl_vfb_0_mem_master_rd_read;          // alt_vip_cl_vfb_0:mem_master_rd_read -> mm_interconnect_0:alt_vip_cl_vfb_0_mem_master_rd_read
	wire         alt_vip_cl_vfb_0_mem_master_rd_readdatavalid; // mm_interconnect_0:alt_vip_cl_vfb_0_mem_master_rd_readdatavalid -> alt_vip_cl_vfb_0:mem_master_rd_readdatavalid
	wire   [6:0] alt_vip_cl_vfb_0_mem_master_rd_burstcount;    // alt_vip_cl_vfb_0:mem_master_rd_burstcount -> mm_interconnect_0:alt_vip_cl_vfb_0_mem_master_rd_burstcount
	wire         alt_vip_cl_vfb_0_mem_master_wr_waitrequest;   // mm_interconnect_0:alt_vip_cl_vfb_0_mem_master_wr_waitrequest -> alt_vip_cl_vfb_0:mem_master_wr_waitrequest
	wire  [31:0] alt_vip_cl_vfb_0_mem_master_wr_address;       // alt_vip_cl_vfb_0:mem_master_wr_address -> mm_interconnect_0:alt_vip_cl_vfb_0_mem_master_wr_address
	wire   [3:0] alt_vip_cl_vfb_0_mem_master_wr_byteenable;    // alt_vip_cl_vfb_0:mem_master_wr_byteenable -> mm_interconnect_0:alt_vip_cl_vfb_0_mem_master_wr_byteenable
	wire         alt_vip_cl_vfb_0_mem_master_wr_write;         // alt_vip_cl_vfb_0:mem_master_wr_write -> mm_interconnect_0:alt_vip_cl_vfb_0_mem_master_wr_write
	wire  [31:0] alt_vip_cl_vfb_0_mem_master_wr_writedata;     // alt_vip_cl_vfb_0:mem_master_wr_writedata -> mm_interconnect_0:alt_vip_cl_vfb_0_mem_master_wr_writedata
	wire   [6:0] alt_vip_cl_vfb_0_mem_master_wr_burstcount;    // alt_vip_cl_vfb_0:mem_master_wr_burstcount -> mm_interconnect_0:alt_vip_cl_vfb_0_mem_master_wr_burstcount
	wire         mm_interconnect_0_sdram_s1_chipselect;        // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;          // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;       // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;           // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;              // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;        // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;     // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;             // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;         // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         rst_controller_reset_out_reset;               // rst_controller:reset_out -> [alt_vip_cl_cps_0:main_reset, alt_vip_cl_crs_0:main_reset, alt_vip_cl_csc_0:main_reset, alt_vip_cl_cvi_0:main_reset_reset, alt_vip_cl_dil_0:av_st_reset, alt_vip_cl_vfb_0:main_reset, alt_vip_cl_vfb_0:mem_reset, alt_vip_clip_1:main_reset, alt_vip_itc_0:rst, alt_vip_scl_0:main_reset, mm_interconnect_0:alt_vip_cl_vfb_0_mem_reset_reset_bridge_in_reset_reset, sdram:reset_n]

	DE10_Standard_VIP_Qsys_alt_vip_cl_cps_0 #(
		.BITS_PER_SYMBOL     (8),
		.USER_PACKET_SUPPORT ("PASSTHROUGH")
	) alt_vip_cl_cps_0 (
		.main_clock           (pll_0_outclk1_clk),                     // main_clock.clk
		.main_reset           (rst_controller_reset_out_reset),        // main_reset.reset
		.din_0_data           (alt_vip_cl_cvi_0_dout_0_data),          //      din_0.data
		.din_0_valid          (alt_vip_cl_cvi_0_dout_0_valid),         //           .valid
		.din_0_startofpacket  (alt_vip_cl_cvi_0_dout_0_startofpacket), //           .startofpacket
		.din_0_endofpacket    (alt_vip_cl_cvi_0_dout_0_endofpacket),   //           .endofpacket
		.din_0_ready          (alt_vip_cl_cvi_0_dout_0_ready),         //           .ready
		.dout_0_data          (alt_vip_cl_cps_0_dout_0_data),          //     dout_0.data
		.dout_0_valid         (alt_vip_cl_cps_0_dout_0_valid),         //           .valid
		.dout_0_startofpacket (alt_vip_cl_cps_0_dout_0_startofpacket), //           .startofpacket
		.dout_0_endofpacket   (alt_vip_cl_cps_0_dout_0_endofpacket),   //           .endofpacket
		.dout_0_ready         (alt_vip_cl_cps_0_dout_0_ready)          //           .ready
	);

	DE10_Standard_VIP_Qsys_alt_vip_cl_crs_0 alt_vip_cl_crs_0 (
		.main_clock         (pll_0_outclk1_clk),                   // main_clock.clk
		.main_reset         (rst_controller_reset_out_reset),      // main_reset.reset
		.din_data           (alt_vip_cl_vfb_0_dout_data),          //        din.data
		.din_valid          (alt_vip_cl_vfb_0_dout_valid),         //           .valid
		.din_startofpacket  (alt_vip_cl_vfb_0_dout_startofpacket), //           .startofpacket
		.din_endofpacket    (alt_vip_cl_vfb_0_dout_endofpacket),   //           .endofpacket
		.din_ready          (alt_vip_cl_vfb_0_dout_ready),         //           .ready
		.dout_data          (alt_vip_cl_crs_0_dout_data),          //       dout.data
		.dout_valid         (alt_vip_cl_crs_0_dout_valid),         //           .valid
		.dout_startofpacket (alt_vip_cl_crs_0_dout_startofpacket), //           .startofpacket
		.dout_endofpacket   (alt_vip_cl_crs_0_dout_endofpacket),   //           .endofpacket
		.dout_ready         (alt_vip_cl_crs_0_dout_ready)          //           .ready
	);

	DE10_Standard_VIP_Qsys_alt_vip_cl_csc_0 alt_vip_cl_csc_0 (
		.main_clock         (pll_0_outclk1_clk),                   // main_clock.clk
		.main_reset         (rst_controller_reset_out_reset),      // main_reset.reset
		.din_data           (alt_vip_cl_crs_0_dout_data),          //        din.data
		.din_valid          (alt_vip_cl_crs_0_dout_valid),         //           .valid
		.din_startofpacket  (alt_vip_cl_crs_0_dout_startofpacket), //           .startofpacket
		.din_endofpacket    (alt_vip_cl_crs_0_dout_endofpacket),   //           .endofpacket
		.din_ready          (alt_vip_cl_crs_0_dout_ready),         //           .ready
		.dout_data          (alt_vip_cl_csc_0_dout_data),          //       dout.data
		.dout_valid         (alt_vip_cl_csc_0_dout_valid),         //           .valid
		.dout_startofpacket (alt_vip_cl_csc_0_dout_startofpacket), //           .startofpacket
		.dout_endofpacket   (alt_vip_cl_csc_0_dout_endofpacket),   //           .endofpacket
		.dout_ready         (alt_vip_cl_csc_0_dout_ready)          //           .ready
	);

	DE10_Standard_VIP_Qsys_alt_vip_cl_cvi_0 #(
		.BPS                           (8),
		.NUMBER_OF_COLOUR_PLANES       (2),
		.COLOUR_PLANES_ARE_IN_PARALLEL (0),
		.SYNC_TO                       (0),
		.MATCH_CTRLDATA_PKT_CLIP_BASIC (0),
		.MATCH_CTRLDATA_PKT_PAD_ADV    (0),
		.OVERFLOW_HANDLING             (0),
		.USE_EMBEDDED_SYNCS            (1),
		.USE_HDMI_DEPRICATION          (0),
		.GENERATE_VID_F                (0),
		.USE_STD                       (0),
		.STD_WIDTH                     (1),
		.GENERATE_ANC                  (0),
		.ANC_DEPTH                     (1),
		.EXTRACT_TOTAL_RESOLUTION      (1),
		.INTERLACED                    (1),
		.H_ACTIVE_PIXELS_F0            (720),
		.V_ACTIVE_LINES_F0             (288),
		.V_ACTIVE_LINES_F1             (288),
		.FIFO_DEPTH                    (2048),
		.CLOCKS_ARE_SAME               (0),
		.USE_CONTROL                   (0)
	) alt_vip_cl_cvi_0 (
		.main_clock_clk                   (pll_0_outclk1_clk),                                 //    main_clock.clk
		.main_reset_reset                 (rst_controller_reset_out_reset),                    //    main_reset.reset
		.dout_0_data                      (alt_vip_cl_cvi_0_dout_0_data),                      //        dout_0.data
		.dout_0_valid                     (alt_vip_cl_cvi_0_dout_0_valid),                     //              .valid
		.dout_0_startofpacket             (alt_vip_cl_cvi_0_dout_0_startofpacket),             //              .startofpacket
		.dout_0_endofpacket               (alt_vip_cl_cvi_0_dout_0_endofpacket),               //              .endofpacket
		.dout_0_ready                     (alt_vip_cl_cvi_0_dout_0_ready),                     //              .ready
		.clocked_video_vid_clk            (alt_vip_cl_cvi_0_clocked_video_vid_clk),            // clocked_video.vid_clk
		.clocked_video_vid_data           (alt_vip_cl_cvi_0_clocked_video_vid_data),           //              .vid_data
		.clocked_video_vid_de             (alt_vip_cl_cvi_0_clocked_video_vid_de),             //              .vid_de
		.clocked_video_vid_datavalid      (alt_vip_cl_cvi_0_clocked_video_vid_datavalid),      //              .vid_datavalid
		.clocked_video_vid_locked         (alt_vip_cl_cvi_0_clocked_video_vid_locked),         //              .vid_locked
		.clocked_video_vid_f              (alt_vip_cl_cvi_0_clocked_video_vid_f),              //              .vid_f
		.clocked_video_vid_v_sync         (alt_vip_cl_cvi_0_clocked_video_vid_v_sync),         //              .vid_v_sync
		.clocked_video_vid_h_sync         (alt_vip_cl_cvi_0_clocked_video_vid_h_sync),         //              .vid_h_sync
		.clocked_video_vid_color_encoding (alt_vip_cl_cvi_0_clocked_video_vid_color_encoding), //              .vid_color_encoding
		.clocked_video_vid_bit_width      (alt_vip_cl_cvi_0_clocked_video_vid_bit_width),      //              .vid_bit_width
		.clocked_video_sof                (alt_vip_cl_cvi_0_clocked_video_sof),                //              .sof
		.clocked_video_sof_locked         (alt_vip_cl_cvi_0_clocked_video_sof_locked),         //              .sof_locked
		.clocked_video_refclk_div         (alt_vip_cl_cvi_0_clocked_video_refclk_div),         //              .refclk_div
		.clocked_video_clipping           (alt_vip_cl_cvi_0_clocked_video_clipping),           //              .clipping
		.clocked_video_padding            (alt_vip_cl_cvi_0_clocked_video_padding),            //              .padding
		.clocked_video_overflow           (alt_vip_cl_cvi_0_clocked_video_overflow)            //              .overflow
	);

	DE10_Standard_VIP_Qsys_alt_vip_cl_dil_0 #(
		.MAX_WIDTH                        (720),
		.MAX_HEIGHT                       (576),
		.USER_PACKET_SUPPORT              ("PASSTHROUGH"),
		.USER_PACKET_FIFO_DEPTH           (0),
		.PIXELS_IN_PARALLEL               (1),
		.BITS_PER_SYMBOL                  (8),
		.NUMBER_OF_COLOR_PLANES           (2),
		.COLOR_PLANES_ARE_IN_PARALLEL     (1),
		.IS_422                           (1),
		.IS_YCBCR                         (1),
		.DEINTERLACE_ALGORITHM            ("BOB"),
		.MOTION_BLEED                     (1),
		.RUNTIME_CONTROL                  (0),
		.MOTION_BPS                       (7),
		.CADENCE_DETECTION                (0),
		.CADENCE_ALGORITHM_NAME           ("CADENCE_32_22_VOF"),
		.CLOCKS_ARE_SEPARATE              (0),
		.MEM_PORT_WIDTH                   (256),
		.WRITE_MASTER_FIFO_DEPTH          (64),
		.WRITE_MASTER_BURST_TARGET        (32),
		.EDI_READ_MASTER_FIFO_DEPTH       (64),
		.EDI_READ_MASTER_BURST_TARGET     (32),
		.MA_READ_MASTER_FIFO_DEPTH        (64),
		.MA_READ_MASTER_BURST_TARGET      (32),
		.MOTION_WRITE_MASTER_FIFO_DEPTH   (64),
		.MOTION_WRITE_MASTER_BURST_TARGET (32),
		.MOTION_READ_MASTER_FIFO_DEPTH    (64),
		.MOTION_READ_MASTER_BURST_TARGET  (32),
		.MEM_BASE_ADDR                    (0)
	) alt_vip_cl_dil_0 (
		.av_st_clock        (pll_0_outclk1_clk),                     // av_st_clock.clk
		.av_st_reset        (rst_controller_reset_out_reset),        // av_st_reset.reset
		.din_data           (alt_vip_cl_cps_0_dout_0_data),          //         din.data
		.din_valid          (alt_vip_cl_cps_0_dout_0_valid),         //            .valid
		.din_startofpacket  (alt_vip_cl_cps_0_dout_0_startofpacket), //            .startofpacket
		.din_endofpacket    (alt_vip_cl_cps_0_dout_0_endofpacket),   //            .endofpacket
		.din_ready          (alt_vip_cl_cps_0_dout_0_ready),         //            .ready
		.dout_data          (alt_vip_cl_dil_0_dout_data),            //        dout.data
		.dout_valid         (alt_vip_cl_dil_0_dout_valid),           //            .valid
		.dout_startofpacket (alt_vip_cl_dil_0_dout_startofpacket),   //            .startofpacket
		.dout_endofpacket   (alt_vip_cl_dil_0_dout_endofpacket),     //            .endofpacket
		.dout_ready         (alt_vip_cl_dil_0_dout_ready)            //            .ready
	);

	DE10_Standard_VIP_Qsys_alt_vip_cl_vfb_0 #(
		.BITS_PER_SYMBOL              (8),
		.NUMBER_OF_COLOR_PLANES       (2),
		.COLOR_PLANES_ARE_IN_PARALLEL (1),
		.PIXELS_IN_PARALLEL           (1),
		.READY_LATENCY                (1),
		.MAX_WIDTH                    (720),
		.MAX_HEIGHT                   (480),
		.CLOCKS_ARE_SEPARATE          (1),
		.MEM_PORT_WIDTH               (32),
		.MEM_BASE_ADDR                (0),
		.BURST_ALIGNMENT              (1),
		.WRITE_FIFO_DEPTH             (512),
		.WRITE_BURST_TARGET           (64),
		.READ_FIFO_DEPTH              (512),
		.READ_BURST_TARGET            (64),
		.WRITER_RUNTIME_CONTROL       (0),
		.READER_RUNTIME_CONTROL       (0),
		.IS_FRAME_WRITER              (0),
		.IS_FRAME_READER              (0),
		.DROP_FRAMES                  (1),
		.REPEAT_FRAMES                (1),
		.DROP_REPEAT_USER             (1),
		.INTERLACED_SUPPORT           (0),
		.CONTROLLED_DROP_REPEAT       (0),
		.DROP_INVALID_FIELDS          (1),
		.MULTI_FRAME_DELAY            (1),
		.IS_SYNC_MASTER               (0),
		.IS_SYNC_SLAVE                (0),
		.USER_PACKETS_MAX_STORAGE     (0),
		.MAX_SYMBOLS_PER_PACKET       (10),
		.NUM_BUFFERS                  (3)
	) alt_vip_cl_vfb_0 (
		.main_clock                  (pll_0_outclk1_clk),                            //    main_clock.clk
		.main_reset                  (rst_controller_reset_out_reset),               //    main_reset.reset
		.mem_clock                   (pll_0_outclk1_clk),                            //     mem_clock.clk
		.mem_reset                   (rst_controller_reset_out_reset),               //     mem_reset.reset
		.din_data                    (alt_vip_clip_1_dout_data),                     //           din.data
		.din_valid                   (alt_vip_clip_1_dout_valid),                    //              .valid
		.din_startofpacket           (alt_vip_clip_1_dout_startofpacket),            //              .startofpacket
		.din_endofpacket             (alt_vip_clip_1_dout_endofpacket),              //              .endofpacket
		.din_ready                   (alt_vip_clip_1_dout_ready),                    //              .ready
		.mem_master_wr_address       (alt_vip_cl_vfb_0_mem_master_wr_address),       // mem_master_wr.address
		.mem_master_wr_burstcount    (alt_vip_cl_vfb_0_mem_master_wr_burstcount),    //              .burstcount
		.mem_master_wr_waitrequest   (alt_vip_cl_vfb_0_mem_master_wr_waitrequest),   //              .waitrequest
		.mem_master_wr_write         (alt_vip_cl_vfb_0_mem_master_wr_write),         //              .write
		.mem_master_wr_writedata     (alt_vip_cl_vfb_0_mem_master_wr_writedata),     //              .writedata
		.mem_master_wr_byteenable    (alt_vip_cl_vfb_0_mem_master_wr_byteenable),    //              .byteenable
		.dout_data                   (alt_vip_cl_vfb_0_dout_data),                   //          dout.data
		.dout_valid                  (alt_vip_cl_vfb_0_dout_valid),                  //              .valid
		.dout_startofpacket          (alt_vip_cl_vfb_0_dout_startofpacket),          //              .startofpacket
		.dout_endofpacket            (alt_vip_cl_vfb_0_dout_endofpacket),            //              .endofpacket
		.dout_ready                  (alt_vip_cl_vfb_0_dout_ready),                  //              .ready
		.mem_master_rd_address       (alt_vip_cl_vfb_0_mem_master_rd_address),       // mem_master_rd.address
		.mem_master_rd_burstcount    (alt_vip_cl_vfb_0_mem_master_rd_burstcount),    //              .burstcount
		.mem_master_rd_waitrequest   (alt_vip_cl_vfb_0_mem_master_rd_waitrequest),   //              .waitrequest
		.mem_master_rd_read          (alt_vip_cl_vfb_0_mem_master_rd_read),          //              .read
		.mem_master_rd_readdata      (alt_vip_cl_vfb_0_mem_master_rd_readdata),      //              .readdata
		.mem_master_rd_readdatavalid (alt_vip_cl_vfb_0_mem_master_rd_readdatavalid)  //              .readdatavalid
	);

	DE10_Standard_VIP_Qsys_alt_vip_clip_1 #(
		.BITS_PER_SYMBOL              (8),
		.NUMBER_OF_COLOR_PLANES       (2),
		.COLOR_PLANES_ARE_IN_PARALLEL (1),
		.PIXELS_IN_PARALLEL           (1),
		.MAX_IN_WIDTH                 (720),
		.MAX_IN_HEIGHT                (576),
		.CLIPPING_METHOD              ("RECTANGLE"),
		.LEFT_OFFSET                  (0),
		.RIGHT_OFFSET                 (10),
		.TOP_OFFSET                   (24),
		.BOTTOM_OFFSET                (10),
		.RECTANGLE_WIDTH              (720),
		.RECTANGLE_HEIGHT             (480),
		.USER_PACKET_SUPPORT          ("PASSTHROUGH"),
		.RUNTIME_CONTROL              (0),
		.LIMITED_READBACK             (0)
	) alt_vip_clip_1 (
		.main_clock         (pll_0_outclk1_clk),                   // main_clock.clk
		.main_reset         (rst_controller_reset_out_reset),      // main_reset.reset
		.din_data           (alt_vip_cl_dil_0_dout_data),          //        din.data
		.din_valid          (alt_vip_cl_dil_0_dout_valid),         //           .valid
		.din_startofpacket  (alt_vip_cl_dil_0_dout_startofpacket), //           .startofpacket
		.din_endofpacket    (alt_vip_cl_dil_0_dout_endofpacket),   //           .endofpacket
		.din_ready          (alt_vip_cl_dil_0_dout_ready),         //           .ready
		.dout_data          (alt_vip_clip_1_dout_data),            //       dout.data
		.dout_valid         (alt_vip_clip_1_dout_valid),           //           .valid
		.dout_startofpacket (alt_vip_clip_1_dout_startofpacket),   //           .startofpacket
		.dout_endofpacket   (alt_vip_clip_1_dout_endofpacket),     //           .endofpacket
		.dout_ready         (alt_vip_clip_1_dout_ready)            //           .ready
	);

	alt_vipitc131_IS2Vid #(
		.NUMBER_OF_COLOUR_PLANES       (3),
		.COLOUR_PLANES_ARE_IN_PARALLEL (1),
		.BPS                           (8),
		.INTERLACED                    (0),
		.H_ACTIVE_PIXELS               (640),
		.V_ACTIVE_LINES                (480),
		.ACCEPT_COLOURS_IN_SEQ         (0),
		.FIFO_DEPTH                    (1280),
		.CLOCKS_ARE_SAME               (0),
		.USE_CONTROL                   (0),
		.NO_OF_MODES                   (1),
		.THRESHOLD                     (639),
		.STD_WIDTH                     (1),
		.GENERATE_SYNC                 (0),
		.USE_EMBEDDED_SYNCS            (0),
		.AP_LINE                       (0),
		.V_BLANK                       (0),
		.H_BLANK                       (0),
		.H_SYNC_LENGTH                 (96),
		.H_FRONT_PORCH                 (16),
		.H_BACK_PORCH                  (48),
		.V_SYNC_LENGTH                 (2),
		.V_FRONT_PORCH                 (10),
		.V_BACK_PORCH                  (33),
		.F_RISING_EDGE                 (0),
		.F_FALLING_EDGE                (0),
		.FIELD0_V_RISING_EDGE          (0),
		.FIELD0_V_BLANK                (0),
		.FIELD0_V_SYNC_LENGTH          (0),
		.FIELD0_V_FRONT_PORCH          (0),
		.FIELD0_V_BACK_PORCH           (0),
		.ANC_LINE                      (0),
		.FIELD0_ANC_LINE               (0)
	) alt_vip_itc_0 (
		.is_clk        (pll_0_outclk1_clk),                         //       is_clk_rst.clk
		.rst           (rst_controller_reset_out_reset),            // is_clk_rst_reset.reset
		.is_data       (alt_vip_scl_0_dout_data),                   //              din.data
		.is_valid      (alt_vip_scl_0_dout_valid),                  //                 .valid
		.is_ready      (alt_vip_scl_0_dout_ready),                  //                 .ready
		.is_sop        (alt_vip_scl_0_dout_startofpacket),          //                 .startofpacket
		.is_eop        (alt_vip_scl_0_dout_endofpacket),            //                 .endofpacket
		.vid_clk       (alt_vip_itc_0_clocked_video_vid_clk),       //    clocked_video.export
		.vid_data      (alt_vip_itc_0_clocked_video_vid_data),      //                 .export
		.underflow     (alt_vip_itc_0_clocked_video_underflow),     //                 .export
		.vid_datavalid (alt_vip_itc_0_clocked_video_vid_datavalid), //                 .export
		.vid_v_sync    (alt_vip_itc_0_clocked_video_vid_v_sync),    //                 .export
		.vid_h_sync    (alt_vip_itc_0_clocked_video_vid_h_sync),    //                 .export
		.vid_f         (alt_vip_itc_0_clocked_video_vid_f),         //                 .export
		.vid_h         (alt_vip_itc_0_clocked_video_vid_h),         //                 .export
		.vid_v         (alt_vip_itc_0_clocked_video_vid_v)          //                 .export
	);

	DE10_Standard_VIP_Qsys_alt_vip_scl_0 alt_vip_scl_0 (
		.main_clock         (pll_0_outclk1_clk),                   // main_clock.clk
		.main_reset         (rst_controller_reset_out_reset),      // main_reset.reset
		.din_data           (alt_vip_cl_csc_0_dout_data),          //        din.data
		.din_valid          (alt_vip_cl_csc_0_dout_valid),         //           .valid
		.din_startofpacket  (alt_vip_cl_csc_0_dout_startofpacket), //           .startofpacket
		.din_endofpacket    (alt_vip_cl_csc_0_dout_endofpacket),   //           .endofpacket
		.din_ready          (alt_vip_cl_csc_0_dout_ready),         //           .ready
		.dout_data          (alt_vip_scl_0_dout_data),             //       dout.data
		.dout_valid         (alt_vip_scl_0_dout_valid),            //           .valid
		.dout_startofpacket (alt_vip_scl_0_dout_startofpacket),    //           .startofpacket
		.dout_endofpacket   (alt_vip_scl_0_dout_endofpacket),      //           .endofpacket
		.dout_ready         (alt_vip_scl_0_dout_ready)             //           .ready
	);

	DE10_Standard_VIP_Qsys_pll_0 pll_0 (
		.refclk   (clk_clk),           //  refclk.clk
		.rst      (~reset_reset_n),    //   reset.reset
		.outclk_0 (clk_sdram_clk),     // outclk0.clk
		.outclk_1 (pll_0_outclk1_clk), // outclk1.clk
		.outclk_2 (clk_vga_clk),       // outclk2.clk
		.outclk_3 (clk_aud_clk),       // outclk3.clk
		.locked   ()                   //  locked.export
	);

	DE10_Standard_VIP_Qsys_sdram sdram (
		.clk            (pll_0_outclk1_clk),                        //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	DE10_Standard_VIP_Qsys_mm_interconnect_0 mm_interconnect_0 (
		.pll_0_outclk1_clk                                      (pll_0_outclk1_clk),                            //                                    pll_0_outclk1.clk
		.alt_vip_cl_vfb_0_mem_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),               // alt_vip_cl_vfb_0_mem_reset_reset_bridge_in_reset.reset
		.alt_vip_cl_vfb_0_mem_master_rd_address                 (alt_vip_cl_vfb_0_mem_master_rd_address),       //                   alt_vip_cl_vfb_0_mem_master_rd.address
		.alt_vip_cl_vfb_0_mem_master_rd_waitrequest             (alt_vip_cl_vfb_0_mem_master_rd_waitrequest),   //                                                 .waitrequest
		.alt_vip_cl_vfb_0_mem_master_rd_burstcount              (alt_vip_cl_vfb_0_mem_master_rd_burstcount),    //                                                 .burstcount
		.alt_vip_cl_vfb_0_mem_master_rd_read                    (alt_vip_cl_vfb_0_mem_master_rd_read),          //                                                 .read
		.alt_vip_cl_vfb_0_mem_master_rd_readdata                (alt_vip_cl_vfb_0_mem_master_rd_readdata),      //                                                 .readdata
		.alt_vip_cl_vfb_0_mem_master_rd_readdatavalid           (alt_vip_cl_vfb_0_mem_master_rd_readdatavalid), //                                                 .readdatavalid
		.alt_vip_cl_vfb_0_mem_master_wr_address                 (alt_vip_cl_vfb_0_mem_master_wr_address),       //                   alt_vip_cl_vfb_0_mem_master_wr.address
		.alt_vip_cl_vfb_0_mem_master_wr_waitrequest             (alt_vip_cl_vfb_0_mem_master_wr_waitrequest),   //                                                 .waitrequest
		.alt_vip_cl_vfb_0_mem_master_wr_burstcount              (alt_vip_cl_vfb_0_mem_master_wr_burstcount),    //                                                 .burstcount
		.alt_vip_cl_vfb_0_mem_master_wr_byteenable              (alt_vip_cl_vfb_0_mem_master_wr_byteenable),    //                                                 .byteenable
		.alt_vip_cl_vfb_0_mem_master_wr_write                   (alt_vip_cl_vfb_0_mem_master_wr_write),         //                                                 .write
		.alt_vip_cl_vfb_0_mem_master_wr_writedata               (alt_vip_cl_vfb_0_mem_master_wr_writedata),     //                                                 .writedata
		.sdram_s1_address                                       (mm_interconnect_0_sdram_s1_address),           //                                         sdram_s1.address
		.sdram_s1_write                                         (mm_interconnect_0_sdram_s1_write),             //                                                 .write
		.sdram_s1_read                                          (mm_interconnect_0_sdram_s1_read),              //                                                 .read
		.sdram_s1_readdata                                      (mm_interconnect_0_sdram_s1_readdata),          //                                                 .readdata
		.sdram_s1_writedata                                     (mm_interconnect_0_sdram_s1_writedata),         //                                                 .writedata
		.sdram_s1_byteenable                                    (mm_interconnect_0_sdram_s1_byteenable),        //                                                 .byteenable
		.sdram_s1_readdatavalid                                 (mm_interconnect_0_sdram_s1_readdatavalid),     //                                                 .readdatavalid
		.sdram_s1_waitrequest                                   (mm_interconnect_0_sdram_s1_waitrequest),       //                                                 .waitrequest
		.sdram_s1_chipselect                                    (mm_interconnect_0_sdram_s1_chipselect)         //                                                 .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (pll_0_outclk1_clk),              //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
